library verilog;
use verilog.vl_types.all;
entity tb_traffic_light is
    generic(
        DURATION        : integer := 1000
    );
end tb_traffic_light;
